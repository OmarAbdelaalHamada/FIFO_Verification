package shared_pkg;
    import FIFO_transaction_pkg::*;
    import FIFO_coverage_pkg::*;
    integer correct_counter = 0;
    integer error_counter   = 0;
    bit test_finished = 0;
endpackage